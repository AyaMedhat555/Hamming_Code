library verilog;
use verilog.vl_types.all;
entity tb_hammingcode is
end tb_hammingcode;
